
architecture ruturt_arc of ruturt is

	signal clock : std_logic;

begin

end ruturt_arc;